
package ConvLoopParam;
    localparam Pix = 3;
    localparam Piy = 3;
    localparam Nif = 2;
    localparam RES = 4;
    localparam kx = 3;
    localparam Pof = 4;
    localparam Tof = 8;
endpackage


package ConvLoopParam;
    localparam Pix = 3;
    localparam Piy = 3;
    localparam Nif = 2;
    localparam RES = 8;
    localparam kx = 3;
endpackage
